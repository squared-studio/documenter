class test_Class#(
    parameter int size = bit [(1):(0)]
);
    function new();

    endfunction
endclass
